-----------------------------------------------------------------------
-- Authors      : Muhammed Tarık YILDIZ <muhammettarikyildiz@gmail.com>
--              : Murat Can Işık <kernet1@hotmail.com>
-- Project      : OSCILLOSCOPE
-- File Name    : signal_process.vhd
-- Title        : Signal Processing
-- Description  :
-----------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY SIGNAL_PROCESS IS

PORT
(
	CLK: IN STD_LOGIC;
	INT1,INT2:IN STD_LOGIC;
	RD1,RD2:OUT STD_LOGIC;
	WR1,WR2:OUT STD_LOGIC;
	ADC_DATA_IN1,ADC_DATA_IN2:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL_RAM_RD_ADDR1: IN STD_LOGIC_VECTOR(11 DOWNTO 0);
	SIGNAL_RAM_RD_DATA1: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL_RAM_RD_ADDR2: IN STD_LOGIC_VECTOR(11 DOWNTO 0);
	SIGNAL_RAM_RD_DATA2: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	VPP_MAX1:OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	VPP_MAX2:OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	VPP_MIN1:OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	VPP_MIN2:OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	PERIODE1:OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	PERIODE2:OUT STD_LOGIC_VECTOR(12 DOWNTO 0)
);
END ENTITY SIGNAL_PROCESS;


ARCHITECTURE ARCH_SIGNAL_PROCESS OF SIGNAL_PROCESS IS
COMPONENT ADC IS

PORT( 
	M_CLK:IN  STD_LOGIC:='0'; 
	INT : IN  STD_LOGIC:='1'; 
	RD  : OUT  STD_LOGIC:='1';
	WR  :OUT STD_LOGIC:='0'; 
	ADC_DATA_IN:IN STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000"; 
	ADC_INT:OUT INTEGER RANGE 0 TO 255;
	ADC_DATA_OUT:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	ADC_ENABLE:OUT STD_LOGIC
	); 

END COMPONENT ADC;

COMPONENT SIGNAL_RAM IS
PORT(	
		CLK: IN STD_LOGIC;
		WRITE_ADRR: IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		READ_ADDR:IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		DATA_IN: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		DATA_OUT:OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		);
END COMPONENT SIGNAL_RAM;
COMPONENT SIGNAL_MEASUREMENT IS 
PORT
(
		CLK: IN STD_LOGIC;
		RST: IN STD_LOGIC;
		ADC_DATA1: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		ADC_DATA2:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		VPPMAX1 : OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
		VPPMAX2 : OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
		VPPMIN1 : OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
		VPPMIN2 : OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
		PERIODE1 : OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
		PERIODE2 : OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
		MAX1_OUT : OUT INTEGER RANGE 0 TO 255;
		MAX2_OUT : OUT INTEGER RANGE 0 TO 255;
		MIN1_OUT : OUT INTEGER RANGE 0 TO 255;
		MIN2_OUT : OUT INTEGER RANGE 0 TO 255
);
END COMPONENT SIGNAL_MEASUREMENT;
SIGNAL WR_ADDR1,WR_ADDR2:STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL DATA_IN1,DATA_IN2:STD_LOGIC_VECTOR(7 DOWNTO 0);

SIGNAL MAX1,MAX2,MIN1,MIN2:INTEGER RANGE 0 TO 255;
SIGNAL ADC_INT1,ADC_INT2:INTEGER RANGE 0 TO 255;
SIGNAL ADC_DATA_OUT1,ADC_DATA_OUT2:STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL ADC_ENABLE1,ADC_ENABLE2:STD_LOGIC;
SIGNAL CNT1,CNT2:INTEGER RANGE 0 TO 4095 := 0;
SIGNAL RST:STD_LOGIC := '0';
SIGNAL COUNT_TIME: INTEGER RANGE 0 TO 50_000_000 := 0;
SIGNAL COUNT_SECOND:INTEGER RANGE 0 TO 3 := 0;
BEGIN
ADC1: ADC PORT MAP(CLK,INT1,RD1,WR1,ADC_DATA_IN1,ADC_INT1,ADC_DATA_OUT1,ADC_ENABLE1);
ADC2: ADC PORT MAP(CLK,INT2,RD2,WR2,ADC_DATA_IN2,ADC_INT2,ADC_DATA_OUT2,ADC_ENABLE2);
SIGNAL_MEASUREMENT_C: SIGNAL_MEASUREMENT PORT MAP(CLK,RST,ADC_DATA_OUT1,ADC_DATA_OUT2,VPP_MAX1,VPP_MAX2,VPP_MIN1,VPP_MIN2,PERIODE1,PERIODE2,MAX1,MAX2,MIN1,MIN2);
SINGAL_RAM1:SIGNAL_RAM PORT MAP(CLK,WR_ADDR1,SIGNAL_RAM_RD_ADDR1,DATA_IN1,SIGNAL_RAM_RD_DATA1);
SIGNAL_RAM2:SIGNAL_RAM PORT MAP(CLK,WR_ADDR2,SIGNAL_RAM_RD_ADDR2,DATA_IN2,SIGNAL_RAM_RD_DATA2);

PROCESS(CLK)
BEGIN
IF RISING_EDGE(CLK) THEN	
	--COUNT TIME
	IF COUNT_TIME = 50_000_000 THEN
		COUNT_TIME <= 0;
		RST <= '1';
	ELSE
		RST <= '0';
		COUNT_TIME <= COUNT_TIME + 1;
	END IF;
	
	IF ADC_ENABLE1 = '1' THEN
		WR_ADDR1 <= STD_LOGIC_VECTOR(TO_UNSIGNED(CNT1,12));
		DATA_IN1 <= ADC_DATA_OUT1;
		IF CNT1 = 4095 AND ADC_INT1-MAX1 < 5 THEN
			CNT1 <= 0;
		ELSIF CNT1 /= 4095 THEN
			CNT1 <= CNT1 + 1;
		END IF;
	END IF;
	
	IF ADC_ENABLE2 = '1' THEN
		WR_ADDR2 <= STD_LOGIC_VECTOR(TO_UNSIGNED(CNT2,12));
		DATA_IN2 <= ADC_DATA_OUT2;
		IF CNT2 = 4095 AND ADC_INT2-MAX2<5 THEN
			CNT2 <= 0;
		ELSIF CNT2 /= 4095  THEN
			CNT2 <= CNT2 + 1;
		END IF;
	END IF;
	
END IF;
END PROCESS;

END ARCHITECTURE ARCH_SIGNAL_PROCESS;