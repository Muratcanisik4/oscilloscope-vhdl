-----------------------------------------------------------------------
-- Authors      : Muhammed Tarık YILDIZ <muhammettarikyildiz@gmail.com>
--              : Murat Can Işık <kernet1@hotmail.com>
-- Project      : OSCILLOSCOPE
-- File Name    : oscilloscope.vhd
-- Title        : Oscilloscope Controller
-- Description  :
------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY OSCILLOSCOPE IS

PORT
(
		CLK:IN STD_LOGIC; -- SYSTEM CLOCK PIN
		INT1,INT2:IN STD_LOGIC; --ADC PINS
		RD1,RD2:OUT STD_LOGIC; -- ADC PINS
		WR1,WR2:OUT STD_LOGIC; -- ADC PINS
		ADC_DATA_IN1:IN STD_LOGIC_VECTOR(7 DOWNTO 0); --ADC PINS
		ADC_DATA_IN2:IN STD_LOGIC_VECTOR(7 DOWNTO 0); --ADC PINS
		VGA_R,VGA_G,VGA_B: OUT STD_LOGIC; -- VGA PINS
		VGA_HSYNC,VGA_VSYNC:OUT STD_LOGIC -- VGA PINS
);

END ENTITY OSCILLOSCOPE;


ARCHITECTURE ARCH_OSCILLOSCOPE OF OSCILLOSCOPE IS
COMPONENT VGA_DRIVER IS
PORT
(
		CLK:IN STD_LOGIC;
		SIGNAL_RAM_ADDR1,SIGNAL_RAM_ADDR2:OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
		SIGNAL_RAM_DATA1,SIGNAL_RAM_DATA2:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		VPPMAX1,VPPMAX2,VPPMIN1,VPPMIN2,PERIODE1,PERIODE2:IN STD_LOGIC_VECTOR(12 DOWNTO 0);
		VGA_R,VGA_G,VGA_B:OUT STD_LOGIC;
		VGA_HSYNC,VGA_VSYNC:OUT STD_LOGIC
);
END COMPONENT VGA_DRIVER;
COMPONENT SIGNAL_PROCESS IS
PORT
(
	CLK: IN STD_LOGIC;
	INT1,INT2:IN STD_LOGIC;
	RD1,RD2:OUT STD_LOGIC;
	WR1,WR2:OUT STD_LOGIC;
	ADC_DATA_IN1,ADC_DATA_IN2:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL_RAM_RD_ADDR1: IN STD_LOGIC_VECTOR(11 DOWNTO 0);
	SIGNAL_RAM_RD_DATA1: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL_RAM_RD_ADDR2: IN STD_LOGIC_VECTOR(11 DOWNTO 0);
	SIGNAL_RAM_RD_DATA2: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	VPP_MAX1:OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	VPP_MAX2:OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	VPP_MIN1:OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	VPP_MIN2:OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	PERIODE1:OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	PERIODE2:OUT STD_LOGIC_VECTOR(12 DOWNTO 0)
);
END COMPONENT SIGNAL_PROCESS;

SIGNAL SIGNAL_RAM_ADDR1,SIGNAL_RAM_ADDR2:STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL SIGNAL_RAM_DATA1,SIGNAL_RAM_DATA2:STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL VPPMAX1,VPPMAX2,VPPMIN1,VPPMIN2,PERIODE1,PERIODE2:STD_LOGIC_VECTOR(12 DOWNTO 0);

BEGIN
VGA_DRIVER_C: VGA_DRIVER PORT MAP(CLK,SIGNAL_RAM_ADDR1,SIGNAL_RAM_ADDR2,SIGNAL_RAM_DATA1,SIGNAL_RAM_DATA2,VPPMAX1,VPPMAX2,VPPMIN1,VPPMIN2,PERIODE1,PERIODE2,VGA_R,VGA_G,VGA_B,VGA_HSYNC,VGA_VSYNC);
SIGNAL_PROCESS_C: SIGNAL_PROCESS PORT MAP(CLK,INT1,INT2,RD1,RD2,WR1,WR2,ADC_DATA_IN1,ADC_DATA_IN2,SIGNAL_RAM_ADDR1,SIGNAL_RAM_DATA1,SIGNAL_RAM_ADDR2,SIGNAL_RAM_DATA2,VPPMAX1,VPPMAX2,VPPMIN1,VPPMIN2,PERIODE1,PERIODE2);
END ARCHITECTURE ARCH_OSCILLOSCOPE;