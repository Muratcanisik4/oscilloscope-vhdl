-----------------------------------------------------------------------
-- Authors      : Muhammed Tarık YILDIZ <muhammettarikyildiz@gmail.com>
--              : Murat Can Işık <kernet1@hotmail.com>
-- Project      : OSCILLOSCOPE
-- File Name    : vga_sync.vhd
-- Title        : VGA Interfacing Unit
-- Description  :
-----------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.std_logic_unsigned.all;
USE IEEE.numeric_std.all;
ENTITY VGA_SYNC IS
PORT(
	CLK: IN STD_LOGIC;
	HSYNC, VSYNC: OUT STD_LOGIC;
	R_OUT, G_OUT, B_OUT: OUT STD_LOGIC;
	R_IN: IN STD_LOGIC;
	G_IN: IN STD_LOGIC;
	B_IN: IN STD_LOGIC;
	PIXEL_H: OUT STD_LOGIC_VECTOR(10 DOWNTO 0);
	PIXEL_V: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
	VPPMIN1,VPPMAX1,VPPMIN2,VPPMAX2: IN STD_LOGIC_VECTOR(12 DOWNTO 0);
	PERIODE1,PERIODE2: IN STD_LOGIC_VECTOR(12 DOWNTO 0)
);
END ENTITY VGA_SYNC;

ARCHITECTURE ARCH_VGA_SYNC OF VGA_SYNC IS

TYPE rom_type_23_126 IS ARRAY (0 TO 2897) OF STD_LOGIC;
SUBTYPE c_array_10_7 IS STD_LOGIC_VECTOR(0 TO 69);-- 10X7
SUBTYPE c_array_5_7 IS STD_LOGIC_VECTOR(0 TO 34);--5X7
SUBTYPE c_array_7_7 IS STD_LOGIC_VECTOR(0 TO 48);--7X7
CONSTANT c_zero: c_array_10_7:=( -- 10x7-
'0','0','0','1','1','1','1','1','0','0',
'0','0','1','1','0','0','0','1','1','0',
'0','1','1','0','0','0','0','0','1','1',
'0','1','1','0','0','0','0','0','1','1',
'0','1','1','0','0','0','0','0','1','1',
'0','0','1','1','0','0','0','1','1','0',
'0','0','0','1','1','1','1','1','0','0');

CONSTANT c_one: c_array_10_7:=( --10x7-
'0','0','0','0','0','1','1','0','0','0',  
'0','0','0','1','1','1','1','0','0','0',
'0','0','0','0','0','1','1','0','0','0',
'0','0','0','0','0','1','1','0','0','0',   
'0','0','0','0','0','1','1','0','0','0',  
'0','0','0','0','0','1','1','0','0','0', 
'0','0','0','1','1','1','1','1','1','0');

CONSTANT c_two: c_array_10_7:=(  --10x7-
'0','0','1','1','1','1','1','1','1','0',
'0','1','1','0','0','0','0','0','1','1',
'0','0','0','0','0','0','0','0','1','1',
'0','0','1','1','1','1','1','1','1','0',
'0','1','1','0','0','0','0','0','0','0',
'0','1','1','0','0','0','0','0','0','0',
'0','1','1','1','1','1','1','1','1','1');

CONSTANT c_three: c_array_10_7:=( --10x7-
'0','0','1','1','1','1','1','1','1','0',
'0','1','1','0','0','0','0','0','1','1',
'0','0','0','0','0','0','0','0','1','1',
'0','0','1','1','1','1','1','1','1','0',
'0','0','0','0','0','0','0','0','1','1',
'0','1','1','0','0','0','0','0','1','1',
'0','0','1','1','1','1','1','1','1','0');

CONSTANT c_four: c_array_10_7:=( --10x7-
'0','1','1','0','0','0','0','0','0','0',
'0','1','1','0','0','0','0','1','1','0',
'0','1','1','0','0','0','0','1','1','0',
'0','1','1','0','0','0','0','1','1','0',
'0','1','1','1','1','1','1','1','1','1',
'0','0','0','0','0','0','0','1','1','0',
'0','0','0','0','0','0','0','1','1','0');

CONSTANT c_five: c_array_10_7:=(--10x7-
'0','1','1','1','1','1','1','1','1','0', 
'0','1','1','0','0','0','0','0','0','0',
'0','1','1','0','0','0','0','0','0','0',
'0','1','1','1','1','1','1','1','0','0', 
'0','0','0','0','0','0','0','1','1','0', 
'0','1','1','0','0','0','0','1','1','0', 
'0','0','1','1','1','1','1','1','0','0'); 

CONSTANT c_six: c_array_10_7:=(--10x7-
'0','0','1','1','1','1','1','1','1','0',
'0','1','1','0','0','0','0','0','1','1',
'0','1','1','0','0','0','0','0','0','0',
'0','1','1','1','1','1','1','1','1','0',
'0','1','1','0','0','0','0','0','1','1',
'0','1','1','0','0','0','0','0','1','1',
'0','0','1','1','1','1','1','1','1','0');

CONSTANT c_seven: c_array_10_7:=( --10x7-
'0','1','1','1','1','1','1','1','1','0', 
'0','1','1','0','0','0','0','1','1','0', 
'0','0','0','0','0','1','1','0','0','0', 
'0','0','0','0','1','1','0','0','0','0', 
'0','0','0','1','1','0','0','0','0','0', 
'0','0','0','1','1','0','0','0','0','0', 
'0','0','0','1','1','0','0','0','0','0'); 

CONSTANT c_eight: c_array_10_7:=( --10x7-
'0','0','1','1','1','1','1','1','1','0',
'0','1','1','0','0','0','0','0','1','1',
'0','1','1','0','0','0','0','0','1','1',
'0','0','1','1','1','1','1','1','1','0',
'0','1','1','0','0','0','0','0','1','1',
'0','1','1','0','0','0','0','0','1','1',
'0','0','1','1','1','1','1','1','1','0');

CONSTANT c_nine: c_array_10_7:=( --10x7-
'0','0','1','1','1','1','1','1','1','0',
'0','1','1','0','0','0','0','0','1','1',
'0','1','1','0','0','0','0','0','1','1',
'0','0','1','1','1','1','1','1','1','1',
'0','0','0','0','0','0','0','0','1','1',
'0','1','1','0','0','0','0','0','1','1',
'0','0','1','1','1','1','1','1','1','0');

CONSTANT c_comma: c_array_5_7:=( --5x7-
'0','0','0','0','0',     
'0','0','0','0','0',     
'0','0','0','0','0',     
'0','1','1','1','1',     
'0','1','1','1','1',     
'0','0','1','1','0',     
'0','1','1','0','0');     

CONSTANT c_m: c_array_10_7:=( --10x7-
'0','0','0','0','0','0','0','0','0','0', 
'0','0','0','0','0','0','0','0','0','0',
'0','1','1','1','1','1','1','1','1','0',
'0','1','1','1','1','1','1','1','1','0',
'0','1','1','1','1','1','1','1','1','0',
'0','1','1','0','1','1','0','1','1','0',
'0','1','1','0','1','1','0','1','1','0'); 
CONSTANT c_u: c_array_10_7:=( --10x7-
'0','0','0','0','0','0','0','0','0','0', 
'0','0','0','0','0','0','0','0','0','0',
'0','1','1','0','0','1','1','0','0','0',
'0','1','1','0','0','1','1','0','0','0',
'0','1','1','0','0','1','1','0','0','0',
'0','1','1','1','1','1','1','0','0','0',
'0','1','1','1','1','1','1','0','0','0'); 

CONSTANT c_plus: c_array_7_7:=( --7x7-
'0','0','0','0','0','0','0',  
'0','0','0','1','1','0','0',   
'0','0','0','1','1','0','0',   
'0','1','1','1','1','1','1',   
'0','0','0','1','1','0','0',   
'0','0','0','1','1','0','0',   
'0','0','0','0','0','0','0'); 

CONSTANT c_minus: c_array_7_7:=( --7x7-
'0','0','0','0','0','0','0', 
'0','0','0','0','0','0','0', 
'0','0','0','0','0','0','0',  
'0','1','1','1','1','1','1',  
'0','0','0','0','0','0','0',  
'0','0','0','0','0','0','0',
'0','0','0','0','0','0','0');  
constant titles:rom_type_23_126:=('0','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','0','1','1','1','1','1','1','1','1','0','0','1','1','1','1','0','0','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','1','1','1','1','1','1','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0',
'0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','1','1','0','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1',
'0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','1','1','0','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0',
'0','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','0','0','0','1','1','1','1','1','1','1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','1','1','0','1','1','1','1','1','1','0','0','0','1','1','0','0','0','0','0','1','1','1','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
'0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','1','1','0','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0',
'0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1',
'0','1','1','0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1','0','1','1','0','0','0','0','0','1','1','0','1','1','1','1','0','0','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0','0','1','1','1','0','0','1','1','1','1','1','1','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0',
'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
'0','1','1','0','0','0','0','0','1','1','0','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','1','0','1','1','0','0','0','0','0','1','1','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1',                                
'0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','1','1','0','1','1','1','0','0','0','1','1','1','0','0','0','1','1','0','1','1','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1',                    
'0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','1','1','0','1','1','1','1','0','1','1','1','1','0','0','1','1','0','0','0','1','1','0','0','0','0','1','1','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1',                                
'0','1','1','0','0','0','0','0','1','1','0','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0','1','1','0','1','1','1','0','1','1','0','1','1','0','0','0','0','0','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',                                 
'0','0','1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','1','1','1','1','1','1','1','1','1','0','0','0','1','1','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1',                               
'0','0','0','1','1','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','1','1','0','0','1','1','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1',                                 
'0','0','0','0','1','1','1','0','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1',                                 
'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
'0','1','1','0','0','0','0','0','1','1','0','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0','1','1','0','0','0','0','0','1','1','0','1','1','1','1','0','1','1','0','0','0','0','1','1','0','0','0','0','0','0','1','1','1','0','1','1','0','0','0','0','0','1','1','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1',                                          
'0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','1','1','0','1','1','1','0','0','0','1','1','1','0','0','1','1','0','0','1','1','1','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1',                                        
'0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','1','1','0','1','1','1','1','0','1','1','1','1','0','0','1','1','0','0','1','1','1','1','0','0','1','1','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1',                                        
'0','1','1','0','0','0','0','0','1','1','0','1','1','1','1','1','1','1','1','0','0','1','1','1','1','1','1','1','1','0','0','1','1','0','1','1','1','0','1','1','0','0','1','1','0','0','1','1','0','1','1','0','1','1','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',                                          
'0','0','1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','1','1','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0',                                        
'0','0','0','1','1','0','1','1','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','1','1','0','0','1','1','0','0','0','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','1',                                          
'0','0','0','0','1','1','1','0','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','1','1','1','1','0','1','1','0','0','0','0','1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0');                                                                                    
SIGNAL HPOS: INTEGER RANGE 0 TO 1040:=0;
SIGNAL VPOS: INTEGER RANGE 0 TO 666:=0;
SIGNAL COUNT_TITLE1: INTEGER RANGE 0 TO 2897 := 0;
SIGNAL COUNT_TITLE2: INTEGER RANGE 0 TO 2897 := 0; 
SIGNAL COUNT: INTEGER RANGE 0 TO 6 := 0;
SUBTYPE LINE_ARRAY IS STD_LOGIC_VECTOR(0 TO 454);
------------------------------------------------------
SIGNAL CHAR_A1:c_array_10_7; -- (+)ABC(K) -- CH1 --PERIODE_TUENCY
SIGNAL CHAR_B1:c_array_10_7;
SIGNAL CHAR_C1:c_array_10_7;
SIGNAL CHAR_MILI_MICRO1: c_array_10_7;
------------------------------------------------------
SIGNAL CHAR_SIGN11:c_array_7_7; -- (+)C,DE --CH1 --VPPMAX
SIGNAL CHAR_C11:c_array_10_7;
SIGNAL CHAR_D11: c_array_10_7;
SIGNAL CHAR_E11: c_array_10_7;
-------------------------------------------------------
SIGNAL CHAR_SIGN12:c_array_7_7; -- (+)C,DE --CH1 --VPPMIN
SIGNAL CHAR_C12:c_array_10_7;
SIGNAL CHAR_D12: c_array_10_7;
SIGNAL CHAR_E12: c_array_10_7;
------------------------------------------------------
SIGNAL CHAR_A2:c_array_10_7; -- (+)ABC(K) -- CH2 --PERIODE_TUENCY
SIGNAL CHAR_B2:c_array_10_7;
SIGNAL CHAR_C2:c_array_10_7;
SIGNAL CHAR_MILI_MICRO2: c_array_10_7;
------------------------------------------------------
SIGNAL CHAR_SIGN21:c_array_7_7; -- (+)C,DE --CH2 --VPPMAX
SIGNAL CHAR_C21:c_array_10_7;
SIGNAL CHAR_D21: c_array_10_7;
SIGNAL CHAR_E21: c_array_10_7;
-------------------------------------------------------
SIGNAL CHAR_SIGN22:c_array_7_7; -- (+)C,DE --CH2 --VPPMIN
SIGNAL CHAR_C22:c_array_10_7;
SIGNAL CHAR_D22: c_array_10_7;
SIGNAL CHAR_E22: c_array_10_7;
---------------------------------------------------------
SIGNAL CHAR_COMMA:c_array_5_7;
---------------------------------------------------------
SIGNAL COUNT_SIGN:INTEGER RANGE 0 TO 48 := 0;
SIGNAL COUNT_A:INTEGER RANGE 0 TO 69 := 0;
SIGNAL COUNT_B:INTEGER RANGE 0 TO 69 := 0;
SIGNAL COUNT_C:INTEGER RANGE 0 TO 69 := 0;
SIGNAL COUNT_COMMA: INTEGER RANGE 0 TO 34 := 0;
SIGNAL COUNT_D: INTEGER RANGE 0 TO 69 := 0;
SIGNAL COUNT_E: INTEGER RANGE 0 TO 69 :=0;
SIGNAL COUNT_KILO: INTEGER RANGE 0 TO 69 := 0;
SHARED VARIABLE R,G,B:STD_LOGIC;
---------------------------------------------------------
FUNCTION CHAR_SELECT (NUMBER : INTEGER RANGE 0 TO 9) RETURN c_array_10_7 IS
BEGIN
	CASE NUMBER IS
		WHEN 0 => RETURN c_zero;
		WHEN 1 => RETURN c_one;
		WHEN 2 => RETURN c_two;
		WHEN 3 => RETURN c_three;
		WHEN 4 => RETURN c_four;
		WHEN 5 => RETURN c_five;
		WHEN 6 => RETURN c_six;
		WHEN 7 => RETURN c_seven;
		WHEN 8 => RETURN c_eight;
		WHEN 9 => RETURN c_nine;
		WHEN OTHERS => NULL;
	END CASE;

END FUNCTION CHAR_SELECT;-- 1(SIGN BIT, 1 NEGATIVE,0 POSITIVE)--VPP 11(LEFT ON THE COMMA)--1111111(RIGHT ON THE COMMA)
--------------------------------------------------------------
PROCEDURE PRINT_SCREEN_VPP(SIGNAL VPP:IN STD_LOGIC_VECTOR(12 DOWNTO 0);SIGNAL C_OUT,D_OUT,E_OUT:OUT c_array_10_7;SIGNAL C_SIGN:OUT c_array_7_7) IS
BEGIN
IF VPP(12) = '1' THEN -- 1 MINUS
	C_SIGN <= c_plus;
	--C_SIGN <= c_minus;
ELSE 
	C_SIGN <= c_plus;
END IF;
C_OUT <= CHAR_SELECT(TO_INTEGER(UNSIGNED(VPP(11 DOWNTO 8))));
D_OUT <= CHAR_SELECT(TO_INTEGER(UNSIGNED(VPP(7 DOWNTO 4))));
E_OUT <= CHAR_SELECT(TO_INTEGER(UNSIGNED(VPP(3 DOWNTO 0))));
END PROCEDURE;
--------------------------------------------------------------
PROCEDURE PRINT_SCREEN_PRIODE(SIGNAL PERIODE_T:IN STD_LOGIC_VECTOR(12 DOWNTO 0);SIGNAL A_OUT,B_OUT,C_OUT,K_OUT:OUT c_array_10_7) IS
VARIABLE COUNT_1,COUNT_2,COUNT_3:INTEGER:= 0;
BEGIN
IF(PERIODE_T(12) = '1') THEN
	K_OUT <= c_m; --ms mili
ELSE
	K_OUT <= c_u; --us micro
END IF;
A_OUT <= CHAR_SELECT(TO_INTEGER(UNSIGNED(PERIODE_T(11 DOWNTO 8)))); 
B_OUT <= CHAR_SELECT(TO_INTEGER(UNSIGNED(PERIODE_T(7 DOWNTO 4))));
C_OUT <= CHAR_SELECT(TO_INTEGER(UNSIGNED(PERIODE_T(3 DOWNTO 0))));
END PROCEDURE;
--------------------------------------------------------------
SIGNAL COUNT_H : STD_LOGIC_VECTOR(10 DOWNTO 0) := "00000000000";
SIGNAL COUNT_V : STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
--------------------------------------------------------------
BEGIN
CHAR_COMMA <= c_comma;
PROCESS(PERIODE1,PERIODE2,VPPMAX1,VPPMIN1,VPPMAX2,VPPMIN2)
BEGIN
PRINT_SCREEN_PRIODE(PERIODE1,CHAR_A1,CHAR_B1,CHAR_C1,CHAR_MILI_MICRO1);
PRINT_SCREEN_PRIODE(PERIODE2,CHAR_A2,CHAR_B2,CHAR_C2,CHAR_MILI_MICRO2);
PRINT_SCREEN_VPP(VPPMAX1,CHAR_C11,CHAR_D11,CHAR_E11,CHAR_SIGN11);
PRINT_SCREEN_VPP(VPPMIN1,CHAR_C12,CHAR_D12,CHAR_E12,CHAR_SIGN12);
PRINT_SCREEN_VPP(VPPMAX2,CHAR_C21,CHAR_D21,CHAR_E21,CHAR_SIGN21);
PRINT_SCREEN_VPP(VPPMIN2,CHAR_C22,CHAR_D22,CHAR_E22,CHAR_SIGN22);
END PROCESS;

PIXEL_H <= COUNT_H;
PIXEL_V <= COUNT_V;

PROCESS(CLK)
VARIABLE ADDR_STD:STD_LOGIC_VECTOR(11 DOWNTO 0) := "000000000000";
VARIABLE HPOS_CLC:INTEGER RANGE 0 TO 360;
BEGIN
	IF (rising_edge(CLK)) THEN
		IF HPOS<=800 AND VPOS<=600 THEN
			IF HPOS >=240 AND HPOS < 600 THEN 
				IF VPOS>66 AND VPOS<=266 THEN --360 X 200 -- CH1 SIGNAL SCREEN
				       R := R_IN;
					   G := '0';
					   B := '0';
				ELSIF VPOS>266 AND VPOS<=466 THEN --360 X 200 -- CH2 SIGNAL SCREEN
					   R := '0';
					   G := '0';
					   B := B_IN;
				ELSE 
					   R := '0';
					   G := '0';
				END IF;
			ELSE
				R:='0';
				G:='0';
				B:='0';
			END IF;
			--INFO PERIODE_TUENCY,VPPMAX,VPPMIN
			IF HPOS>=600 AND HPOS<=725 AND VPOS<=266 AND VPOS>=244 THEN
				R:= TITLES(COUNT_TITLE1);
				G:= '0';
				B:= '0';
				IF COUNT_TITLE1 = 2897 THEN
					COUNT_TITLE1 <= 0;
				ELSE
					COUNT_TITLE1 <= COUNT_TITLE1 + 1;
				END IF;
			ELSIF HPOS>=600 AND HPOS<=725 AND VPOS<=466 AND VPOS>=444 THEN
				R:='0';
				G:='0';
				B:=TITLES(COUNT_TITLE2);
				IF COUNT_TITLE2 = 2897 THEN
					COUNT_TITLE2 <= 0;
				ELSE
					COUNT_TITLE2 <= COUNT_TITLE2 + 1;
				END IF;
			ELSIF HPOS > 725 AND HPOS <= 790 THEN
				    IF VPOS<=266 AND VPOS>=244 THEN -- CHANNEL 1
						IF VPOS<=250 AND VPOS>=244 THEN -- PERIODE_TUENCY
							IF HPOS>=726  AND HPOS<=735 THEN --CHAR_A
								R := CHAR_A1(COUNT_A);
								G := '0';
								B := '0';
								IF COUNT_A = 69 THEN
									COUNT_A <= 0;
								ELSE
									COUNT_A <= COUNT_A + 1;
								END IF;
							ELSIF HPOS>=736 AND HPOS <=745 THEN --CHAR_B
								R := CHAR_B1(COUNT_B);
								G := '0';
								B := '0';
								IF COUNT_B = 69 THEN
									COUNT_B <= 0;
								ELSE
									COUNT_B <= COUNT_B + 1;
								END IF;
							ELSIF HPOS>=746 AND HPOS<=755 THEN -- CHAR C
								R := CHAR_C1(COUNT_C);
								G := '0';
								B := '0';
								IF COUNT_C = 69 THEN
									COUNT_C <= 0;
								ELSE
									COUNT_C <= COUNT_C + 1;
								END IF;
							ELSIF HPOS>=756 AND HPOS<=765 THEN --CHAR KILO
								R := CHAR_MILI_MICRO1(COUNT_KILO);
								G := '0';
								B := '0';
								IF COUNT_KILO = 69 THEN
									COUNT_KILO <= 0;
								ELSE
									COUNT_KILO <= COUNT_KILO + 1;
								END IF;
							END IF;
						ELSIF VPOS<=258 AND VPOS>=252 THEN -- VPPMAX
							IF HPOS>=726  AND HPOS<=732 THEN --CHAR_SIGN
								R := CHAR_SIGN11(COUNT_SIGN);
								G := '0';
								B := '0';
								IF COUNT_SIGN = 48 THEN
									COUNT_SIGN <= 0;
								ELSE
									COUNT_SIGN <= COUNT_SIGN + 1;
								END IF;
							
							ELSIF HPOS>=733 AND HPOS<=742 THEN -- CHAR C
								R := CHAR_C11(COUNT_C);
								G := '0';
								B := '0';
								IF COUNT_C = 69 THEN
									COUNT_C <= 0;
								ELSE
									COUNT_C <= COUNT_C + 1;
								END IF;
							ELSIF HPOS>=743 AND HPOS<=747 THEN --CHAR COMMA
								R := CHAR_COMMA(COUNT_COMMA);
								G := '0';
								B := '0';
								IF COUNT_COMMA = 34 THEN
									COUNT_COMMA <= 0;
								ELSE
									COUNT_COMMA <= COUNT_COMMA + 1;
								END IF;
							ELSIF HPOS>=748 AND HPOS<=757 THEN --CHAR D
								R := CHAR_D11(COUNT_D);
								G := '0';
								B := '0';
								IF COUNT_D = 69 THEN
									COUNT_D <= 0;
								ELSE
									COUNT_D <= COUNT_D + 1;
								END IF;
							ELSIF HPOS>=758 AND HPOS<=767 THEN --CHAR E
								R := CHAR_E11(COUNT_E);
								G := '0';
								B := '0';
								IF COUNT_E = 69 THEN
									COUNT_E <= 0;
								ELSE
									COUNT_E <= COUNT_E + 1;
								END IF;
							ELSE
								R:='0';
								G:='0';
								B:='0';
							END IF;
						ELSIF VPOS<=266 AND VPOS>=260 THEN -- VPPMIN
							IF HPOS>=726  AND HPOS<=732 THEN --CHAR_SIGN
								R := CHAR_SIGN12(COUNT_SIGN);
								G := '0';
								b := '0';
								IF COUNT_SIGN = 48 THEN
									COUNT_SIGN <= 0;
								ELSE
									COUNT_SIGN <= COUNT_SIGN + 1;
								END IF;
							
							ELSIF HPOS>=733 AND HPOS<=742 THEN -- CHAR C
								R := CHAR_C12(COUNT_C);
								G := '0';
								b := '0';
								IF COUNT_C = 69 THEN
									COUNT_C <= 0;
								ELSE
									COUNT_C <= COUNT_C + 1;
								END IF;
							ELSIF HPOS>=743 AND HPOS<=747 THEN --CHAR COMMA
								R := CHAR_COMMA(COUNT_COMMA);
								G := '0';
								b := '0';
								IF COUNT_COMMA = 34 THEN
									COUNT_COMMA <= 0;
								ELSE
									COUNT_COMMA <= COUNT_COMMA + 1;
								END IF;
							ELSIF HPOS>=748 AND HPOS<=757 THEN --CHAR D
								R := CHAR_D12(COUNT_D);
								G := '0';
								b := '0';
								IF COUNT_D = 69 THEN
									COUNT_D <= 0;
								ELSE
									COUNT_D <= COUNT_D + 1;
								END IF;
							ELSIF HPOS>=758 AND HPOS<=767 THEN --CHAR E
								R := CHAR_E12(COUNT_E);
								G := '0';
								b := '0';
								IF COUNT_E = 69 THEN
									COUNT_E <= 0;
								ELSE
									COUNT_E <= COUNT_E + 1;
								END IF;
							ELSE
								R:='0';
								G:='0';
								B:='0';
							END IF;
						END IF;
				    ELSIF VPOS<=466 AND VPOS>=444 THEN -- CHANNEL 2
						IF VPOS<=450 AND VPOS>=444 THEN -- PERIODE_TUENCY
							IF HPOS>=726  AND HPOS<=735 THEN --CHAR_A
								B := CHAR_A2(COUNT_A);
								G := '0';
								R := '0';
								IF COUNT_A = 69 THEN
									COUNT_A <= 0;
								ELSE
									COUNT_A <= COUNT_A + 1;
								END IF;
							ELSIF HPOS>=736 AND HPOS <=745 THEN --CHAR_B
								B := CHAR_B2(COUNT_B);
								G := '0';
								R := '0';
								IF COUNT_B = 69 THEN
									COUNT_B <= 0;
								ELSE
									COUNT_B <= COUNT_B + 1;
								END IF;
							ELSIF HPOS>=746 AND HPOS<=755 THEN -- CHAR C
								B := CHAR_C2(COUNT_C);
								G := '0';
								R := '0';
								IF COUNT_C = 69 THEN
									COUNT_C <= 0;
								ELSE
									COUNT_C <= COUNT_C + 1;
								END IF;
							ELSIF HPOS>=756 AND HPOS<=765 THEN --CHAR KILO
								B := CHAR_MILI_MICRO2(COUNT_KILO);
								G := '0';
								R := '0';
								IF COUNT_KILO = 69 THEN
									COUNT_KILO <= 0;
								ELSE
									COUNT_KILO <= COUNT_KILO + 1;
								END IF;
							END IF;
						ELSIF VPOS<=458 AND VPOS>=452 THEN -- VPPMAX
							IF HPOS>=726  AND HPOS<=732 THEN --CHAR_SIGN
								B := CHAR_SIGN21(COUNT_SIGN);
								G := '0';
								R := '0';
								IF COUNT_SIGN = 48 THEN
									COUNT_SIGN <= 0;
								ELSE
									COUNT_SIGN <= COUNT_SIGN + 1;
								END IF;

							ELSIF HPOS>=733 AND HPOS<=742 THEN -- CHAR C
								B := CHAR_C21(COUNT_C);
								G := '0';
								R := '0';
								IF COUNT_C = 69 THEN
									COUNT_C <= 0;
								ELSE
									COUNT_C <= COUNT_C + 1;
								END IF;
							ELSIF HPOS>=743 AND HPOS<=747 THEN --CHAR COMMA
								B := CHAR_COMMA(COUNT_COMMA);
								G := '0';
								R := '0';
								IF COUNT_COMMA = 34 THEN
									COUNT_COMMA <= 0;
								ELSE
									COUNT_COMMA <= COUNT_COMMA + 1;
								END IF;
							ELSIF HPOS>=748 AND HPOS<=757 THEN --CHAR D
								B := CHAR_D21(COUNT_D);
								G := '0';
								R := '0';
								IF COUNT_D = 69 THEN
									COUNT_D <= 0;
								ELSE
									COUNT_D <= COUNT_D + 1;
								END IF;
							ELSIF HPOS>=758 AND HPOS<=767 THEN --CHAR E
								B := CHAR_E21(COUNT_E);
								G := '0';
								R := '0';
								IF COUNT_E = 69 THEN
									COUNT_E <= 0;
								ELSE
									COUNT_E <= COUNT_E + 1;
								END IF;
							ELSE
								R:='0';
								G:='0';
								B:='0';
							END IF;
						ELSIF VPOS<=466 AND VPOS>=460 THEN -- VPPMIN
							IF HPOS>=726  AND HPOS<=732 THEN --CHAR_SIGN
								B := CHAR_SIGN22(COUNT_SIGN);
								G := '0';
								R := '0';
								IF COUNT_SIGN = 48 THEN
									COUNT_SIGN <= 0;
								ELSE
									COUNT_SIGN <= COUNT_SIGN + 1;
								END IF;
							
							ELSIF HPOS>=733 AND HPOS<=742 THEN -- CHAR C
								B := CHAR_C22(COUNT_C);
								G := '0';
								R := '0';
								IF COUNT_C = 69 THEN
									COUNT_C <= 0;
								ELSE
									COUNT_C <= COUNT_C + 1;
								END IF;
							ELSIF HPOS>=743 AND HPOS<=747 THEN --CHAR COMMA
								B := CHAR_COMMA(COUNT_COMMA);
								G := '0';
								R := '0';
								IF COUNT_COMMA = 34 THEN
									COUNT_COMMA <= 0;
								ELSE
									COUNT_COMMA <= COUNT_COMMA + 1;
								END IF;
							ELSIF HPOS>=748 AND HPOS<=757 THEN --CHAR D
								B := CHAR_D22(COUNT_D);
								G := '0';
								R := '0';
								IF COUNT_D = 69 THEN
									COUNT_D <= 0;
								ELSE
									COUNT_D <= COUNT_D + 1;
								END IF;
							ELSIF HPOS>=758 AND HPOS<=767 THEN --CHAR E
								B := CHAR_E22(COUNT_E);
								G := '0';
								R := '0';
								IF COUNT_E = 69 THEN
									COUNT_E <= 0;
								ELSE
									COUNT_E <= COUNT_E + 1;
								END IF;
							ELSE
								R:='0';
								G:='0';
								B:='0';
							END IF;
						END IF;
					ELSE
						-- R:='0';
						-- G:='0';
						-- B:='0';
					END IF;
			END IF;
		END IF;
		IF (HPOS<1040) THEN
			HPOS<=HPOS+1;
			COUNT_H <= COUNT_H + '1';
		ELSE
			HPOS<=0;
			COUNT_H <= "00000000000";
			IF (VPOS<666) THEN
				VPOS<=VPOS+1;
				COUNT_V <= COUNT_V + '1';
			ELSE
				VPOS<=0;
				COUNT_V <= "0000000000";
			END IF;
		END IF;
 
		IF (HPOS>56 AND HPOS<176) THEN
			HSYNC<='0';
		ELSE	
			HSYNC<='1';
		END IF;
 
		IF (VPOS>0 AND VPOS<43) THEN -- maybe 37>x<43
			VSYNC<='0';
		ELSE	
			VSYNC<='1';
		END IF;
		IF ((HPOS>0 AND HPOS<240) OR (VPOS>0 AND VPOS<66)) THEN
			R:='0';
			G:='0';
			B:='0';
		END IF;
	END IF;
	R_OUT <= R;
	G_OUT <= G;
	B_OUT <= B;
END PROCESS;
END ARCHITECTURE ARCH_VGA_SYNC;